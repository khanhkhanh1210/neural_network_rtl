module neuron(
	input logic [7:0] x,w_in
	input clk,w_en
	output logic [7:0] w_out
);
rom weight_value(1'b1,w_in,clk,w_en,
always@(posedge clk) begin
	
always@*
	
