module testop();
reg [3:0] a_i,b_i;
wire [3:0] sum_o;
reg c_in;
wire c_out;
endmodule
